

module PYTEST(
    inout  wire b,
    inout  wire d,
    inout  wire g,
    inout  wire s
);

endmodule
